// adder 


module adder 
